// ============================================================================
// top_module
// ----------------------------------------------------------------------------
// Description:
//   Connects the AXI Read Address/Data channels to the reordering logic,
//   utilizing FIFOs to decouple the flow stages and an allocator for unique IDs.
//
// Component Flow:
// 1. AXI Master (axi_ar_in) -> incoming_request_fifo
// 2. incoming_request_fifo -> ar_id_ordering_unit (gets UID from allocator)
// 3. ar_id_ordering_unit -> outgoing_request_fifo
// 4. outgoing_request_fifo -> AXI Slave (axi_ar_out)
//
// 5. AXI Slave (axi_r_in) -> incoming_response_fifo
// 6. incoming_response_fifo -> r_id_ordering_unit (stores in response_park/WM)
// 7. r_id_ordering_unit -> outgoing_response_fifo (releases ordered data)
// 8. outgoing_response_fifo -> AXI Master (axi_r_out)
//
// Allocator (allocator_tag_map) is shared by ar_id_ordering_unit (alloc) and
// r_id_ordering_unit (free + restored ID lookup).

//TODO: match all r_if and ar_if
//TODO: implement everything marked as TODO in the code below
//TODO: count how many cycles it takes for a request to go from axi_ar_in to axi_ar_out
//TODO: count how many cycles it takes for a response to go from axi_r_in to axi_r_out
//TODO: check if r_id_ordering_unit needs FSM like ar_id_ordering_unit
//TODO: add the "last" signal to response_park and every where it's missing and check what happens with multi-beat requests/responses
// ============================================================================
module top_module #(
    parameter int ID_WIDTH          = 4,
    parameter int DATA_WIDTH        = 64,
    parameter int RESP_WIDTH        = 2,
    parameter int TAG_WIDTH         = 4,  // Internal tag width
    parameter int MAX_OUTSTANDING   = 16, // Must match sub-modules
    parameter int ADDR_WIDTH        = 32,
    parameter int LEN_WIDTH         = 8
)(
    input  logic clk,
    input  logic rst,

    // AXI Read Address Channel (AR) Master Interface (Input to this module)
    ar_if.receiver axi_ar_in, //TODO: need to add more fields according to Gil's slides or AXI protocol document
    ar_if.sender    axi_ar_out,

    // AXI Read Data Channel (R) Slave Interface (Output from this module)
    r_if.sender     axi_r_out, //TODO: need to add more fields according to Gil's slides or AXI protocol document
    r_if.receiver   axi_r_in 
);

    // ------------------------------------------------------------------------
    // Derived Parameters
    // ------------------------------------------------------------------------
    localparam int NUM_ROWS = $bits(MAX_OUTSTANDING);
    localparam int NUM_COLS = $bits(MAX_OUTSTANDING);
    localparam int ROW_W = $bits(NUM_ROWS);
    localparam int COL_W = $bits(NUM_COLS);
    localparam int UID_W = ROW_W + COL_W; // Unique ID width

    // Define AXI Read Address fields structure for FIFOs
    // This combines the fields passed from axi_ar_in to axi_ar_out
    typedef struct packed {
        logic [ID_WIDTH-1:0]  id;
        logic [ADDR_WIDTH-1:0] addr;
        logic [LEN_WIDTH-1:0]  len;
        logic [2:0]            size;
        logic [1:0]            burst;
        // NOTE: Add ARQOS/ARCACHE/etc. fields here if needed by ar_if
    } axi_ar_fields_t;

    // Define AXI Read Data fields structure for FIFOs
    // This is the struct of the usual metadata, minus 'valid' and 'ready'
    typedef struct packed {
        logic [ID_WIDTH-1:0] id;
        logic [DATA_WIDTH-1:0] data;
        logic [RESP_WIDTH-1:0] resp;
        logic last;
        logic [TAG_WIDTH-1:0] tagid;
    } axi_r_payload_t;


    // ------------------------------------------------------------------------
    // Allocator Signals (Used by allocator_tag_map, ar_id_ordering_unit, r_id_ordering_unit)
    // ------------------------------------------------------------------------
    logic                 alloc_req;         // from AR unit
    logic [ID_WIDTH-1:0]  alloc_in_id;       // from AR unit
    logic                 alloc_gnt;         // to AR unit
    logic [UID_W-1:0]     alloc_unique_id;   // to AR unit
    logic                 tag_map_full;      // to incoming_request_fifo (TODO: Implement in allocator_tag_map)

    logic                 free_req;          // from R unit
    logic [UID_W-1:0]     free_unique_id;    // from R unit
    logic [ID_WIDTH-1:0]  restored_id;       // to R unit
    logic                 free_ack;

    // ------------------------------------------------------------------------
    // AR Request FIFO Interfaces (axi_ar_fields_t payload)
    // ------------------------------------------------------------------------

    // FIFO 1: Incoming Request FIFO
    axi_ar_fields_t fifo1_in_data;
    logic fifo1_in_valid;
    logic fifo1_in_ready; // Backpressure to axi_ar_in
    axi_ar_fields_t fifo1_out_data;
    logic fifo1_out_valid; // Input to ar_id_ordering_unit
    logic fifo1_out_ready; // From ar_id_ordering_unit
    logic fifo1_full;      // Backpressure to axi_ar_in

    // FIFO 2: Outgoing Request FIFO
    axi_ar_fields_t fifo2_in_data; // From ar_id_ordering_unit
    logic fifo2_in_valid;  // From ar_id_ordering_unit
    logic fifo2_in_ready;  // Backpressure to ar_id_ordering_unit
    axi_ar_fields_t fifo2_out_data;
    logic fifo2_out_valid; // Input to axi_ar_out
    logic fifo2_out_ready; // From axi_ar_out

    // ------------------------------------------------------------------------
    // R Response FIFO Interfaces (axi_r_payload_t payload)
    // ------------------------------------------------------------------------

    // FIFO 3: Incoming Response FIFO
    axi_r_payload_t fifo3_in_data;
    logic fifo3_in_valid;
    logic fifo3_in_ready; // Backpressure to axi_r_in
    axi_r_payload_t fifo3_out_data; // Input to r_id_ordering_unit
    logic fifo3_out_valid;          // Input to r_id_ordering_unit
    logic fifo3_out_ready;          // From r_id_ordering_unit
    logic fifo3_full;               // Backpressure to axi_r_in

    // FIFO 4: Outgoing Response FIFO
    axi_r_payload_t fifo4_in_data;  // From r_id_ordering_unit
    logic fifo4_in_valid;           // From r_id_ordering_unit
    logic fifo4_in_ready;           // Backpressure to r_id_ordering_unit
    axi_r_payload_t fifo4_out_data;
    logic fifo4_out_valid;          // Input to axi_r_out
    logic fifo4_out_ready;          // From axi_r_out

    // ------------------------------------------------------------------------
    // r_id_ordering_unit and response_park Signals
    // ------------------------------------------------------------------------
    logic                 wm_write_en;
    logic [UID_W-1:0]     wm_write_uid;
    axi_r_payload_t       wm_write_payload; // Payload to response_park

    logic                 wm_release_en;
    logic [UID_W-1:0]     wm_release_uid;
    logic                 wm_release_gnt;   // From response_park
    axi_r_payload_t       wm_release_payload; // Data from response_park
    
    logic                 r_park_full; // Backpressure to incoming_response_fifo (TODO: Implement in response_park)


    // ========================================================================
    // AXI to FIFO and FIFO to AXI Connections
    // ========================================================================

    // --- AXI AR Input to FIFO 1 ---
    assign axi_ar_in.ready  = fifo1_in_ready; // Backpressure from FIFO 1

    assign fifo1_in_valid   = axi_ar_in.valid;
    assign fifo1_in_data.id = axi_ar_in.id;
    assign fifo1_in_data.addr = axi_ar_in.addr;
    assign fifo1_in_data.len = axi_ar_in.len;
    assign fifo1_in_data.size = axi_ar_in.size;
    assign fifo1_in_data.burst = axi_ar_in.burst;

    // --- FIFO 2 to AXI AR Output ---
    assign fifo2_out_ready  = axi_ar_out.ready; // Backpressure to FIFO 2

    assign axi_ar_out.valid = fifo2_out_valid;
    assign axi_ar_out.id    = fifo2_out_data.id; // UID
    assign axi_ar_out.addr  = fifo2_out_data.addr;
    assign axi_ar_out.len   = fifo2_out_data.len;
    assign axi_ar_out.size  = fifo2_out_data.size;
    assign axi_ar_out.burst = fifo2_out_data.burst;


    // --- AXI R Input to FIFO 3 ---
    assign axi_r_in.ready   = fifo3_in_ready; // Backpressure from FIFO 3

    // Note: r_if struct contains fields matching axi_r_payload_t
    assign fifo3_in_valid   = axi_r_in.valid;
    assign fifo3_in_data.id    = axi_r_in.id; // This is the UID
    assign fifo3_in_data.data  = axi_r_in.data;
    assign fifo3_in_data.resp  = axi_r_in.resp;
    assign fifo3_in_data.last  = axi_r_in.last;
    assign fifo3_in_data.tagid = axi_r_in.tagid;

    // --- FIFO 4 to AXI R Output ---
    assign fifo4_out_ready  = axi_r_out.ready; // Backpressure to FIFO 4

    assign axi_r_out.valid  = fifo4_out_valid;
    assign axi_r_out.id     = fifo4_out_data.id; // This is the original ID
    assign axi_r_out.data   = fifo4_out_data.data;
    assign axi_r_out.resp   = fifo4_out_data.resp;
    assign axi_r_out.last   = fifo4_out_data.last;
    assign axi_r_out.tagid  = fifo4_out_data.tagid; // The internal tag ID is passed through


    // ========================================================================
    // 1. allocator_tag_map Instantiation
    // ========================================================================
    allocator #(
        .ID_WIDTH(ID_WIDTH),
        .MAX_OUTSTANDING(MAX_OUTSTANDING)
    ) i_allocator_tag_map (
        .clk             (clk),
        .rst             (rst),
        .alloc_req       (alloc_req),
        .in_orig_id           (alloc_in_id),
        .alloc_gnt       (alloc_gnt),
        .unique_id       (alloc_unique_id),
        .id_matrix_full    (tag_map_full), // TODO: allocator_tag_map.sv needs to implement this signal
        .free_req        (free_req),
        .unique_id_to_free (free_unique_id),
        .restored_id     (restored_id),
        .free_ack        (free_ack)
    );

    // ========================================================================
    // 2. ar_id_ordering_unit Instantiation
    // ========================================================================
    // Takes request from FIFO 1, requests UID, and pushes translated request to FIFO 2
    ar_id_ordering_unit #(
        .ID_WIDTH  (ID_WIDTH),
        .UID_WIDTH (UID_W),
        .ADDR_WIDTH(ADDR_WIDTH),
        .LEN_WIDTH (LEN_WIDTH)
    ) i_ar_id_ordering_unit (
        .clk             (clk),
        .rst             (rst),

        // AXI AR from FIFO 1 (input master side)
        .s_ar.valid      (fifo1_out_valid),
        .s_ar.ready      (fifo1_out_ready),
        .s_ar.id         (fifo1_out_data.id),
        .s_ar.addr       (fifo1_out_data.addr),
        .s_ar.len        (fifo1_out_data.len),
        .s_ar.size       (fifo1_out_data.size),
        .s_ar.burst      (fifo1_out_data.burst),

        // AXI AR to FIFO 2 (output slave side - UID is the ID)
        .m_ar.valid      (fifo2_in_valid),
        .m_ar.ready      (fifo2_in_ready),
        .m_ar.id         (fifo2_in_data.id),      // Unique ID output
        .m_ar.addr       (fifo2_in_data.addr),
        .m_ar.len        (fifo2_in_data.len),
        .m_ar.size       (fifo2_in_data.size),
        .m_ar.burst      (fifo2_in_data.burst),

        // Allocator interface
        .alloc_req       (alloc_req),
        .alloc_in_id     (alloc_in_id),
        .alloc_gnt       (alloc_gnt),
        .unique_id       (alloc_unique_id)
    );
    // Note: The ar_id_ordering_unit is designed to take the request directly
    // and not from a FIFO, so we treat the FIFO output handshake as the
    // master side handshake (s_ar.valid/ready). 
    //TODO: change that, ar_id_ordering_unit should not behave like master

    // ========================================================================
    // 3. r_response_waiting_memory (response_park) Instantiation
    // ========================================================================
    // Stores out-of-order responses until requested by r_id_ordering_unit
    response_park #(
        .NUM_ROWS       (NUM_ROWS),
        .NUM_COLS       (NUM_COLS),
        .MAX_REQ        (MAX_OUTSTANDING),
        .DATA_WIDTH     (DATA_WIDTH),
        .RESP_WIDTH     (RESP_WIDTH),
        .ID_WIDTH       (ID_WIDTH),
        .TAG_WIDTH      (TAG_WIDTH)
    ) i_r_response_waiting_memory (
        .clk            (clk),
        .rst            (rst),
        // ENQUEUE (from r_id_ordering_unit when OOO)
        .in_valid       (wm_write_en),
        .in_ready       (/* r_park_full is used to determine readiness */), // Unused in this direction
                                                                            //TODO: delete this signal from response_park.sv
        .in_uid         (wm_write_uid),
        .in_data        (wm_write_payload.data),
        .in_resp        (wm_write_payload.resp),
        .in_orig_id     (wm_write_payload.id),
        .in_tagid       (wm_write_payload.tagid),
        // ALLOCATE (from r_id_ordering_unit to release ordered data)
        .alloc_req      (wm_release_en),
        .alloc_uid      (wm_release_uid),
        // FREE (r_id_ordering_unit/allocator takes care of free)
        .free_req       (free_req),
        .id_to_release  (free_unique_id),
        // OUTPUT
        .alloc_gnt      (wm_release_gnt),
        .out_data       (wm_release_payload.data),
        .out_resp       (wm_release_payload.resp),
        .out_orig_id    (wm_release_payload.id),
        .out_tagid      (wm_release_payload.tagid),
        // Ack/Status
        .free_ack       (/* unused */), //TODO: figure out if needed
        // TODO: needed 'not full' signal from response_park
        // I will use an internal signal from response_park for backpressure.
        .full           (r_park_full) // Assume response_park has a 'full' output
    );

    // ========================================================================
    // 4. r_id_ordering_unit Instantiation
    // ========================================================================
    // Takes response from FIFO 3, reorders, and pushes ordered response to FIFO 4
    r_id_ordering_unit #(
        .ID_WIDTH         (ID_WIDTH),
        .MAX_OUTSTANDING  (MAX_OUTSTANDING),
        .NUM_ROWS         (NUM_ROWS),
        .NUM_COLS         (NUM_COLS),
        .UID_W            (UID_W)
    ) i_r_id_ordering_unit (
        .clk             (clk),
        .rst             (rst),

        // Incoming response (from FIFO 3)
        .resp_valid      (fifo3_out_valid),
        .r_in.ready      (fifo3_out_ready),
        .resp_uid        (fifo3_out_data.id), // UID
        .r_in.id         (fifo3_out_data.id),
        .r_in.data       (fifo3_out_data.data),
        .r_in.resp       (fifo3_out_data.resp),
        .r_in.last       (fifo3_out_data.last),
        .r_in.tagid      (fifo3_out_data.tagid),

        // Outgoing response (to FIFO 4)
        .release_valid   (fifo4_in_valid),
        .r_out.ready     (fifo4_in_ready),
        .r_out.id        (fifo4_in_data.id),  // Original ID output
        .r_out.data      (fifo4_in_data.data),
        .r_out.resp      (fifo4_in_data.resp),
        .r_out.last      (fifo4_in_data.last),
        .r_out.tagid     (fifo4_in_data.tagid),

        // Allocator/Free interface (needs restored_id from allocator_tag_map)
        .restored_id     (restored_id), // TODO: r_id_ordering_unit.sv needs this input to set r_out.id. add this unput signal to r_id_ordering_unit.sv

        // Waiting memory interface (to/from response_park)
        .wm_write_en     (wm_write_en),
        .wm_write_uid    (wm_write_uid),
        // wm_write_data is the data that is being passed to the waiting memory.
        // The r_id_ordering_unit instantiates an r_if.sender for this.
        .wm_write_data.valid (wm_write_payload.valid), // Connect valid/data from r_id_ordering_unit to response_park
        .wm_write_data.id    (wm_write_payload.id),
        .wm_write_data.data  (wm_write_payload.data),
        .wm_write_data.resp  (wm_write_payload.resp),
        .wm_write_data.last  (wm_write_payload.last),
        .wm_write_data.tagid (wm_write_payload.tagid),

        .wm_release_en   (wm_release_en),
        .wm_release_uid  (wm_release_uid),
        // wm_release_data is the data returned from the waiting memory.
        // The r_id_ordering_unit instantiates an r_if.receiver for this.
        .wm_release_data.valid (wm_release_gnt),  // wm_release_data.valid is effectively alloc_gnt from response_park
        .wm_release_data.id    (wm_release_payload.id),
        .wm_release_data.data  (wm_release_payload.data),
        .wm_release_data.resp  (wm_release_payload.resp),
        .wm_release_data.last  (1'b1), // response_park doesn't have 'last', assume 1 beat response for simplicity //TODO: add last to everything
        .wm_release_data.tagid (wm_release_payload.tagid),

        // Backpressure from response_park
        .wm_full         (r_park_full), // Backpressure from response_park.sv. TODO: r_id_ordering_unit.sv needs this input.

        // Free request to allocator
        .free_req        (free_req),
        .free_uid        (free_unique_id)
    );

    // Explicitly connect r_id_ordering_unit's payload to wm_write_payload
    // The r_id_ordering_unit uses r_if.sender for wm_write_data,
    // which has its own logic/data signals, so we need to bridge them.
    // However, the r_id_ordering_unit.sv is designed to drive the signals
    // directly. We must adjust the connection to match the response_park input.
    // The current r_id_ordering_unit code drives the wm_write_data signals
    // on its output modport, which needs to be captured here and passed to
    // response_park's 'in' signals.

    assign wm_write_payload.id    = i_r_id_ordering_unit.wm_write_data.id;
    assign wm_write_payload.data  = i_r_id_ordering_unit.wm_write_data.data;
    assign wm_write_payload.resp  = i_r_id_ordering_unit.wm_write_data.resp;
    assign wm_write_payload.last  = i_r_id_ordering_unit.wm_write_data.last;
    assign wm_write_payload.tagid = i_r_id_ordering_unit.wm_write_data.tagid;
    assign wm_write_payload.valid = i_r_id_ordering_unit.wm_write_data.valid;
    
    // Explicitly connect r_id_ordering_unit's release input from wm_release_payload
    // The r_id_ordering_unit uses r_if.receiver for wm_release_data,
    // which is essentially the output of response_park (alloc_gnt/out_*)

    // Note: the r_id_ordering_unit assumes its r_if.receiver output 'ready'
    // is wired back to response_park, but response_park uses a request/grant pulse.
    // We assume the r_id_ordering_unit does not need to backpressure the response_park
    // and simply consumes the data when 'wm_release_en' and 'wm_release_gnt' are both high.
    //TODO: perhaps change signals accordingly in r_id_ordering_unit.sv and response_park.sv


    // ========================================================================
    // 5. FIFO Instantiations (Using Generic Placeholder)
    // ========================================================================

    // FIFO 1: incoming_request_fifo (AXI AR fields)
    // Push condition: axi_ar_in.valid & ~fifo1_full (implied by fifo1_in_ready)
    // Pop condition: allocator_tag_map is not full (implied by ~tag_map_full)
    // suggestion: implement with standard fifo. below that is a non-standard fifo control.
    // Standard FIFO: Push when in_valid & in_ready. Pop when out_valid & out_ready.
    // We override the push/pop readiness logic below.
    fifo_module #(.D_WIDTH($bits(axi_ar_fields_t)), .DEPTH(16)) i_fifo_ar_in (
        .clk        (clk),
        .rst        (rst),
        .data_in    (fifo1_in_data),
        .valid_in   (fifo1_in_valid),
        .ready_out  (fifo1_in_ready), // Backpressure to axi_ar_in
        .data_out   (fifo1_out_data),
        .valid_out  (fifo1_out_valid),
        .ready_in   (fifo1_out_ready), // Backpressure from ar_id_ordering_unit
        .full       (fifo1_full),
        .empty      (/* unused */)
    );

    // FIFO 2: outgoing_request_fifo (AXI AR fields with UID)
    // Push condition: ar_id_ordering_unit is ready (implied by fifo2_in_ready)
    // Pop condition: axi_ar_out.ready is high
    fifo_module #(.D_WIDTH($bits(axi_ar_fields_t)), .DEPTH(16)) i_fifo_ar_out (
        .clk        (clk),
        .rst        (rst),
        .data_in    (fifo2_in_data),
        .valid_in   (fifo2_in_valid),
        .ready_out  (fifo2_in_ready), // Backpressure to ar_id_ordering_unit
        .data_out   (fifo2_out_data),
        .valid_out  (fifo2_out_valid),
        .ready_in   (fifo2_out_ready), // Pop condition: axi_ar_out.ready
        .full       (/* unused */),
        .empty      (/* unused */)
    );

    // FIFO 3: incoming_response_fifo (AXI R payload)
    // Push condition: axi_r_in.valid & ~fifo3_full (implied by fifo3_in_ready)
    // Pop condition: response can be consumed by r_id_ordering_unit
    fifo_module #(.D_WIDTH($bits(axi_r_payload_t)), .DEPTH(16)) i_fifo_r_in (
        .clk        (clk),
        .rst        (rst),
        .data_in    (fifo3_in_data),
        .valid_in   (fifo3_in_valid),
        .ready_out  (fifo3_in_ready), // Backpressure to axi_r_in
        .data_out   (fifo3_out_data),
        .valid_out  (fifo3_out_valid),
        .ready_in   (fifo3_out_ready), // Pop condition: r_id_ordering_unit consumption
        .full       (fifo3_full),
        .empty      (/* unused */)
    );

    // FIFO 4: outgoing_response_fifo (AXI R payload - original ID)
    // Push condition: r_id_ordering_unit releases a response
    // Pop condition: axi_r_out.ready is high
    fifo_module #(.D_WIDTH($bits(axi_r_payload_t)), .DEPTH(16)) i_fifo_r_out (
        .clk        (clk),
        .rst        (rst),
        .data_in    (fifo4_in_data),
        .valid_in   (fifo4_in_valid),
        .ready_out  (fifo4_in_ready), // Backpressure to r_id_ordering_unit
        .data_out   (fifo4_out_data),
        .valid_out  (fifo4_out_valid),
        .ready_in   (fifo4_out_ready), // Pop condition: axi_r_out.ready
        .full       (/* unused */),
        .empty      (/* unused */)
    );

    // ========================================================================
    // Custom FIFO Flow Control Logic (Overrides Standard Pop/Push)
    // ========================================================================

    // FIFO 1 Pop Control: Pop request when ar_id_ordering_unit is ready (fifo1_out_ready is high)
    // AND the allocator is not full. The ar_id_ordering_unit is a single-entry
    // pipeline that requests the UID, so it becomes ready when it can accept a
    // new request AND the allocator can grant it (preventing deadlock by
    // only accepting if a UID can be granted).
    // The ar_id_ordering_unit handles its own backpressure (s_ar.ready).
    // TODO: We need a check for allocator_tag_map not full (~tag_map_full)
    // to be part of the pop condition for FIFO 1.
    // The current ar_id_ordering_unit has its own backpressure logic (s_ar.ready).
    // For now, we connect FIFO 1 output ready to ar_id_ordering_unit input ready.
    // A more complex implementation would involve checking tag_map_full here
    // or allowing ar_id_ordering_unit to check it before asserting ready.
    // Given the current ar_id_ordering_unit, the backpressure is internal to it.
    // We assume ar_id_ordering_unit ready signal (fifo1_out_ready) implicitly includes
    // the tag map fullness check to prevent deadlock.
    // If our intent is to connect tag_map_full to the FIFO, we must:
    // assign fifo1_out_ready = i_ar_id_ordering_unit.s_ar.ready & ~tag_map_full;
    // but the ar_id_ordering_unit does not expose a ready signal for S_AR.
    // Therefore, we trust the ar_id_ordering_unit's internal logic for now.
    // We will use the output ready signal of the ar_id_ordering_unit.

    // The ar_id_ordering_unit is meant to accept the AR fields directly.
    // We treat its s_ar.ready as the FIFO's pop ready signal.
    assign fifo1_out_ready = i_ar_id_ordering_unit.s_ar.ready;

    // FIFO 3 Pop Control: Pop response when r_id_ordering_unit can consume it.
    // The r_id_ordering_unit accepts a response if:
    // 1. It's a direct hit (and can be immediately released to FIFO 4)
    // 2. It's an out-of-order miss, AND the response_park (wm) is not full.
    // TODO: We need pop if (hit in r_id_ordering_unit) OR (response_park not full).
    // The r_id_ordering_unit.sv does not expose an explicit ready signal for its input.
    // We assume the internal logic of r_id_ordering_unit implicitly drives
    // the ready signal high when it is ready to consume (based on the FIFO pop conditions).
    // We assume a ready signal will be implemented in r_id_ordering_unit.
    // For now, we create a placeholder signal that would be the output ready:
    logic r_id_ordering_unit_ready; // This signal must be driven by r_id_ordering_unit
    assign fifo3_out_ready = r_id_ordering_unit_ready;
    
    // We must pass the necessary information to r_id_ordering_unit so it can drive its ready.
    // The current r_id_ordering_unit does not have a ready input/output.
    // The connection is currently: r_in.ready (from r_id_ordering_unit) -> fifo3_out_ready
    // Since r_if is a receiver modport:
    // assign fifo3_out_ready = i_r_id_ordering_unit.r_in.ready; // The r_if receiver modport for r_in has an output ready.

    // Let's rely on the definition in r_id_ordering_unit.sv:
    // .r_in, r_if.receiver
    // The r_if receiver modport has an output 'ready'.
    assign fifo3_out_ready = i_r_id_ordering_unit.r_in.ready; // The 'ready' signal from r_if.receiver modport is an output.


endmodule
